/*
write_back.sv
This module implements the mux for the write back stage. 
*/

module write_back
    (
        input wire [31:0] pc_result,
        input wire [31:0] alu_result,
        input wire [31:0] data_result,
        input wire [1:0] source_select,
        output logic [31:0] write_result
    );

// Local Parameters
localparam ALU      = 0;
localparam PC       = 2;
localparam D_Mem    = 3;

always_comb
begin
    casex(source_select)
        ALU: write_result = alu_result;
        PC: write_result = pc_result;
        D_Mem: write_result = data_result;
        default: write_result = alu_result;
    endcase
end

endmodule