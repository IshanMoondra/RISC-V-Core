`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06.11.2023 10:47:44
// Design Name: 
// Module Name: rv32_registers
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
//This Module defines the 32 Registers present in the RV32I instruction set. 
//This Module does not have the Program Counter. 
//The Program Counter Module will be defined seperately.

//Probably needs RF Bypass: Added 29th Dec 2024

module rv32_register_file
    (
        input clk,
        input rst_n,
        // input pc_halt,
        input write_reg,
        input [4:0] sel_s1,
        input [4:0] sel_s2,
        input [4:0] sel_d1,
        input wire [31:0] reg_d1,
        output logic [31:0] reg_s1,
        output logic [31:0] reg_s2
    );

// Thirty Two 32bit Registers for RV32 ISA requirement    
reg [31:0] registers [0:31];
logic [5:0] count;
logic [31:0] rf_s1; 
logic [31:0] rf_s2;

// Changing to synchronous negative edge triggered reset
// to facilitate BRAM implementation in Artix 7 FPGAs
// always@(posedge clk, negedge rst_n)
always@(posedge clk)
begin    
    if (!rst_n)
        begin
            rf_s1 <= 0;
            rf_s2 <= 0;
            // Setting $Zero to 0. Doesn't work??
            // registers[0] <= 0;
            // Better way to reset the entire RF without wasting the count variable?
            for (count = 0; count < 32; count = count + 1)
                registers[count] <= 0;
        end
    else
        begin
            // Registered Outputs
            rf_s1 <= (sel_s1 == 0) ? (0) : (registers[sel_s1]);
            rf_s2 <= (sel_s2 == 0) ? (0) : (registers[sel_s2]);            
            // Moving the write condition to negedge clock.  
        end            
end

always @( negedge clk )
begin : RF_Write
    // Register File Input
    // Conditionally Writing to Register File based on write_reg signal
    // Also checking if Destination is not $0. 
    if (write_reg && (sel_d1 != 0))
        registers[sel_d1] <= reg_d1;    
end

// Register File Outputs with RF Bypass
// Note if Synopsys removes $Zero Register or not.
assign reg_s1 = (write_reg && (sel_s1 == sel_d1)) ? reg_d1 : rf_s1;
assign reg_s2 = (write_reg && (sel_s2 == sel_d1)) ? reg_d1 : rf_s2;

endmodule
